module clock_gen(clock);       //module name
input clock;                   // port declaration
endmodule
